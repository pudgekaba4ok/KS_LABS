// Arithmetic-Logic Block (ALB) with specified micro-operations
module alb (
    input wire clk,              // Clock for input registers
    input wire reset,            // Synchronous reset
    input wire [3:0] R_in,       // Input operand R
    input wire [3:0] S_in,       // Input operand S
    input wire CI,               // Carry-in
    input wire [1:0] I,          // Control input (I4, I3)
    output reg [3:0] F_ALB,      // Result output
    output wire CO,              // Carry out
    output wire VO,              // Overflow
    output wire NO,              // Negative flag
    output wire ZO               // Zero flag
);

    // Input buffer registers
    reg [3:0] R_reg, S_reg;
    reg CI_reg;
    reg [1:0] I_reg;

    // Internal signals for operations
    wire [3:0] sum_result, sub_result, or_result, and_not_result;
    wire sum_co, sub_co, sum_vo, sub_vo;

    // Input registers
    always @(posedge clk or posedge reset) begin
        if (reset) begin
            R_reg <= 4'b0;
            S_reg <= 4'b0;
            CI_reg <= 1'b0;
            I_reg <= 2'b0;
        end else begin
            R_reg <= R_in;
            S_reg <= S_in;
            CI_reg <= CI;
            I_reg <= I;
        end
    end

    // Arithmetic operations
    assign {sum_co, sum_result} = R_reg + S_reg + CI_reg;
    assign {sub_co, sub_result} = R_reg - S_reg - 1 + CI_reg;

    // Logical operations
    assign or_result       = R_reg | S_reg;
    assign and_not_result  = (~R_reg) & S_reg;

    // Overflow calculation
    assign sum_vo = (R_reg[3] == S_reg[3]) && (sum_result[3] != R_reg[3]);
    assign sub_vo = (R_reg[3] != S_reg[3]) && (sub_result[3] != R_reg[3]);

    // Result multiplexer
    always @(*) begin
        case (I_reg)
            2'b00: F_ALB = or_result;
            2'b01: F_ALB = sum_result;
            2'b10: F_ALB = and_not_result;
            2'b11: F_ALB = sub_result;
            default: F_ALB = 4'b0000;
        endcase
    end

    // Flag generation
    assign CO = (I_reg == 2'b01) ? sum_co :
            (I_reg == 2'b11) ? ~sub_co : 1'b0;

    assign VO = (I_reg == 2'b01) ? sum_vo :
                (I_reg == 2'b11) ? sub_vo : 1'b0;

    assign NO = F_ALB[3];             // Negative flag (MSB)
    assign ZO = (F_ALB == 4'b0000);   // Zero flag

endmodule
