library verilog;
use verilog.vl_types.all;
entity test_sum is
end test_sum;
