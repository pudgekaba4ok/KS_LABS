library verilog;
use verilog.vl_types.all;
entity tb_sum_7r is
end tb_sum_7r;
