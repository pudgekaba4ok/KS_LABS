library verilog;
use verilog.vl_types.all;
entity tb_multiplex8_1 is
end tb_multiplex8_1;
