module reference_model (
    input [3:0] R,
    input [3:0] S,
    input CI,
    input [1:0] I,
    output reg [3:0] ref_F_ALB,
    output reg ref_CO,
    output reg ref_VO,
    output reg ref_NO,
    output reg ref_ZO
);

    reg [4:0] temp;

    always @(*) begin
        case (I)
            2'b00: begin // R ? S
                ref_F_ALB = R | S;
                ref_CO = 0;
                ref_VO = 0;
            end
            2'b01: begin // R + S + CI
                temp = R + S + CI;
                ref_F_ALB = temp[3:0];
                ref_CO = temp[4];
                ref_VO = (R[3] == S[3]) && (ref_F_ALB[3] != R[3]);
            end
            2'b10: begin // �R & S
                ref_F_ALB = (~R) & S;
                ref_CO = 0;
                ref_VO = 0;
            end
            2'b11: begin // R - S - 1 + CI
                temp = R - S - 1 + CI;
                ref_F_ALB = temp[3:0];
                ref_CO = ~temp[4];  
                ref_VO = (R[3] != S[3]) && (ref_F_ALB[3] != R[3]);
            end
            default: begin
                ref_F_ALB = 4'b0000;
                ref_CO = 0;
                ref_VO = 0;
            end
        endcase
        ref_NO = ref_F_ALB[3];
        ref_ZO = (ref_F_ALB == 4'b0000);
    end

endmodule