library verilog;
use verilog.vl_types.all;
entity alb_tb is
end alb_tb;
